module ROM
	(
		input [31:0] Address_in,
		output reg [31:0] Instruction
	);

	always@(*)
	begin 
		case (Address_in)
			0: Instruction = 32'b10000000000000010000011000001010;//-- Addi r1 ,r0 ,1546
			4: Instruction = 32'b00000100000000010001000000000000;//-- Add  r2 ,r0 ,r1
			8: Instruction = 32'b00001100000000010001100000000000;//-- sub r3 ,r0 ,r1
			12: Instruction = 32'b00010100010000110010000000000000;//-- And r4 ,r2 ,r3
			16: Instruction = 32'b10000100011001010001101000110100;//-- Subi r5 ,r3 ,6708
			20: Instruction = 32'b00011000011001000010100000000000;//-- or r5 ,r3 ,r4
			24: Instruction = 32'b00011100101000000011000000000000;//-- nor  r6 ,r5 ,r0
			28: Instruction = 32'b00011100100000000101100000000000;//-- nor  r11 ,r4 ,r0
			32: Instruction = 32'b00001100101001010010100000000000;//-- sub r5 ,r5 ,r5
			36: Instruction = 32'b10000000000000010000010000000000;//-- Addi  r1 ,r0 ,1024
			40: Instruction = 32'b10010100001000100000000000000000;//-- st r2 ,r1 ,0
			44: Instruction = 32'b10010000001001010000000000000000;//-- ld r5 ,r1 ,0
			48: Instruction = 32'b10100000101000000000000000000001;//-- Bez r5 ,1
			52: Instruction = 32'b00100000101000010011100000000000;//-- xor r7 ,r5 ,r1
			56: Instruction = 32'b00100000101000010000000000000000;//-- xor r0 ,r5 ,r1
			60: Instruction = 32'b00100100011010110011100000000000;//-- sla r7 ,r3 ,r11
			64: Instruction = 32'b00101000011010110100000000000000;//-- sll r8 ,r3 ,r11
			68: Instruction = 32'b00101100011001000100100000000000;//-- sra r9 ,r3 ,r4
			72: Instruction = 32'b00110000011001000101000000000000;//-- srl r10 ,r3 ,r4
			76: Instruction = 32'b10010100001000110000000000000100;//-- st r3 ,r1 ,4
			80: Instruction = 32'b10010100001001000000000000001000;//-- st r4 ,r1 ,8
			84: Instruction = 32'b10010100001001010000000000001100;//-- st r5 ,r1 ,12
			88: Instruction = 32'b10010100001001100000000000010000;//-- st r6 ,r1 ,16
			92: Instruction = 32'b10010000001010110000000000000100;//-- ld r11 ,r1 ,4
			96: Instruction = 32'b10010100001001110000000000010100;//-- st r7 ,r1 ,20
			100: Instruction = 32'b10010100001010000000000000011000;//-- st r8 ,r1 ,24
			104: Instruction = 32'b10010100001010010000000000011100;//-- st r9 ,r1 ,28
			108: Instruction = 32'b10010100001010100000000000100000;//-- st r10 ,r1 ,32
			112: Instruction = 32'b10010100001010110000000000100100;//-- st r11 ,r1 ,36
			116: Instruction = 32'b10000000000000010000000000000011;//-- Addi  r1 ,r0 ,3
			120: Instruction = 32'b10000000000001000000010000000000;//-- Addi r4 ,r0 ,1024
			124: Instruction = 32'b10000000000000100000000000000000;//-- Addi  r2 ,r0 ,0
			128: Instruction = 32'b10000000000000110000000000000001;//-- Addi  r3 ,r0 ,1
			132: Instruction = 32'b10000000000010010000000000000010;//-- Addi  r9 ,r0 ,2
			136: Instruction = 32'b00101000011010010100000000000000;//-- sll r8 ,r3 ,r9
			140: Instruction = 32'b00000100100010000100000000000000;//-- Add  r8 ,r4 ,r8
			144: Instruction = 32'b10010001000001010000000000000000;//-- ld r5 ,r8 ,0
			148: Instruction = 32'b10010001000001101111111111111100;//-- ld r6 ,r8 ,-4
			152: Instruction = 32'b00001100101001100100100000000000;//-- sub  r9 ,r5 ,r6
			156: Instruction = 32'b10000000000010101000000000000000;//-- Addi  r10 ,r0 ,0x8000
			160: Instruction = 32'b10000000000010110000000000010000;//-- Addi r11 ,r0 ,16
			164: Instruction = 32'b00101001010010110101000000000000;//-- sll r10 ,r1 ,r11
			168: Instruction = 32'b00010101001010100100100000000000;//-- And  r9 ,r9 ,r10
			172: Instruction = 32'b10100001001000000000000000000010;//-- Bez r9 ,2
			176: Instruction = 32'b10010101000001011111111111111100;//-- st r5 ,r8 ,-4
			180: Instruction = 32'b10010101000001100000000000000000;//-- st r6 ,r8 ,0
			184: Instruction = 32'b10000000011000110000000000000001;//-- Addi  r3 ,r3 ,1
			188: Instruction = 32'b10100100001000111111111111110001;//-- BNE r1 ,r3 ,-15
			192: Instruction = 32'b10000000010000100000000000000001;//-- Addi  r2 ,r2 ,1
			196: Instruction = 32'b10100100001000101111111111101110;//-- BNE r1 ,r2 ,-18
			200: Instruction = 32'b10000000000000010000010000000000;//-- Addi  r1 ,r0 ,1024
			204: Instruction = 32'b10010000001000100000000000000000;//-- ld ,r2 ,r1 ,0
			208: Instruction = 32'b10010000001000110000000000000100;//-- ld ,r3 ,r1 ,4
			212: Instruction = 32'b10010000001001000000000000001000;//-- ld ,r4 ,r1 ,8
			216: Instruction = 32'b10010000001001000000001000001000;//-- ld ,r4 ,r1 ,520
			220: Instruction = 32'b10010000001001000000010000001000;//-- ld ,r4 ,r1 ,1023
			224: Instruction = 32'b10010000001001010000000000001100;//-- ld ,r5 ,r1 ,12
			228: Instruction = 32'b10010000001001100000000000010000;//-- ld ,r6 ,r1 ,16
			232: Instruction = 32'b10010000001001110000000000010100;//-- ld ,r7 ,r1 ,20
			236: Instruction = 32'b10010000001010000000000000011000;//-- ld ,r8 ,r1 ,24
			240: Instruction = 32'b10010000001010010000000000011100;//-- ld ,r9 ,r1 ,28
			244: Instruction = 32'b10010000001010100000000000100000;//-- ld ,r10,r1 ,32
			248: Instruction = 32'b10010000001010110000000000100100;//-- ld ,r11,r1 ,36
			252: Instruction = 32'b10101000000000001111111111111111;//-- JMP  -1
		endcase
	end

endmodule // ROM